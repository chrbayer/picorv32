/*
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 */

`ifdef PICOSOC_V
`error "artya7c.v must be read before picosoc.v!"
`endif

module artya7c (
	input clk,

	output ser_tx,
	input ser_rx,

	output [7:0] leds,

	output flash_csb,
	output flash_clk,
	inout  [3:0] flash_io
);
	reg vio_reset = 1'b0;

	parameter unsigned VIO_WIDTH = 8;
	wire [VIO_WIDTH-1:0] vio_in;
	wire [VIO_WIDTH-1:0] vio_out;

	vio vio (
		.clk (clk),
		.probe_in0 (vio_in),
		.probe_out0 (vio_out));

	parameter unsigned ILA_WIDTH = 32;
	wire [ILA_WIDTH-1:0] ila_in;

	assign ila_in[0] = resetn;
	assign ila_in[1] = vio_reset;
	assign ila_in[2] = ser_rx;
	assign ila_in[3] = ser_tx;

	assign ila_in[8-1:4] = flash_io_do;
	assign ila_in[12-1:8] = flash_io_oe;
	assign ila_in[16-1:12] = flash_io_di;

	assign ila_in[16] = flash_csb;
	assign ila_in[17] = flash_clk;

	ila ila (
		.clk (clk),
		.probe0 (ila_in));

	assign vio_in = leds;
	always @(posedge clk) vio_reset <= vio_out[0];

	reg [13:0] reset_cnt = 0;
	wire resetn = &reset_cnt & !vio_reset;

	always @(posedge clk) begin
		reset_cnt <= reset_cnt + !resetn;
	end

	wire [3:0] flash_io_oe, flash_io_do, flash_io_di;

	genvar i;
	for (i=0; i<4; i=i+1) begin
		assign flash_io_di[i] = flash_io[i];
		assign flash_io[i] = flash_io_oe[i] ? flash_io_do[i] : 1'bZ;
	end

	wire        iomem_valid;
	reg         iomem_ready;
	wire [3:0]  iomem_wstrb;
	wire [31:0] iomem_addr;
	wire [31:0] iomem_wdata;
	reg  [31:0] iomem_rdata;

	reg [31:0] gpio;
	assign leds = gpio[7:0];

	always @(posedge clk) begin
		if (!resetn) begin
			gpio <= 0;
		end else begin
			iomem_ready <= 0;
			if (iomem_valid && !iomem_ready && iomem_addr[31:24] == 8'h 03) begin
				iomem_ready <= 1;
				iomem_rdata <= gpio;
				if (iomem_wstrb[0]) gpio[ 7: 0] <= iomem_wdata[ 7: 0];
				if (iomem_wstrb[1]) gpio[15: 8] <= iomem_wdata[15: 8];
				if (iomem_wstrb[2]) gpio[23:16] <= iomem_wdata[23:16];
				if (iomem_wstrb[3]) gpio[31:24] <= iomem_wdata[31:24];
			end
		end
	end

	wire flash_io0_oe, flash_io0_do, flash_io0_di;
	wire flash_io1_oe, flash_io1_do, flash_io1_di;
	wire flash_io2_oe, flash_io2_do, flash_io2_di;
	wire flash_io3_oe, flash_io3_do, flash_io3_di;

	assign flash_io_oe = {flash_io3_oe, flash_io2_oe, flash_io1_oe, flash_io0_oe};
	assign flash_io_do = {flash_io3_do, flash_io2_do, flash_io1_do, flash_io0_do};
	assign {flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di} = flash_io_di;
	
	parameter integer MEM_WORDS = 256;

	picosoc #(
		.BARREL_SHIFTER(0),
		.ENABLE_MULDIV(0),
		.MEM_WORDS(MEM_WORDS)
	) soc (
		.clk          (clk         ),
		.resetn       (resetn      ),

		.ser_tx       (ser_tx      ),
		.ser_rx       (ser_rx      ),

		.flash_csb    (flash_csb   ),
		.flash_clk    (flash_clk   ),

		.flash_io0_oe (flash_io0_oe),
		.flash_io1_oe (flash_io1_oe),
		.flash_io2_oe (flash_io2_oe),
		.flash_io3_oe (flash_io3_oe),

		.flash_io0_do (flash_io0_do),
		.flash_io1_do (flash_io1_do),
		.flash_io2_do (flash_io2_do),
		.flash_io3_do (flash_io3_do),

		.flash_io0_di (flash_io0_di),
		.flash_io1_di (flash_io1_di),
		.flash_io2_di (flash_io2_di),
		.flash_io3_di (flash_io3_di),

		.irq_5        (1'b0        ),
		.irq_6        (1'b0        ),
		.irq_7        (1'b0        ),

		.iomem_valid  (iomem_valid ),
		.iomem_ready  (iomem_ready ),
		.iomem_wstrb  (iomem_wstrb ),
		.iomem_addr   (iomem_addr  ),
		.iomem_wdata  (iomem_wdata ),
		.iomem_rdata  (iomem_rdata )
	);
endmodule
